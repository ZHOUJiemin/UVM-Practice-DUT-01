//Testbench Top
//Description: UVM practice on DUT 01
//Modification History
//Date          Author          Description
//2015.12.22    ZHOU Jiemin     First created

//Source Code Starts Here------------------------------------
module tb_top();

  //interface instantiation

  //dut instantiation

  //test instantiation

  //config database

  //run test
  
endmodule
